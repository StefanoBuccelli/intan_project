`timescale 1ns/1ps

module TB_cust_comp();
 
    localparam header_magic_number=64'h0F0E0D0C0B0A09080706050403020100;
 
    reg         clk=0;
    reg         reset = 0;
    reg         data_write;
    reg  [15:0] data_to_write;
    wire [15:0] data_out;
    wire        data_out_valid;
    wire [ 7:0] trig_stim;
    wire        computing;
    reg  [15:0] pipein;
    reg         pipein_en;
    reg         pipeout_en;
    wire [15:0] pipeout;
    reg  [15:0] cfg=16'h0000;
    reg  [ 7:0] stream_en;
    wire [15:0] status;
 
 
    CUST_ARCH  #(
        .BOARD_ID                  (16'h0123),
        .BOARD_VERSION             (16'h4567), 
        .HEADER_MAGIC_NUMBER       (header_magic_number)
        )
    custom_proc_architecture
        (
        .clk                       (clk),
        .reset                     (reset),
        .FIFO_write_to             (data_write),         
        .FIFO_data_in              (data_to_write),
        .comp_data_out_valid       (data_out_valid),       
        .comp_data_out             (data_out),         
        .trig_stim                 (trig_stim),             
        .computing                 (computing),     
        .pipe_in_data              (pipein),      
        .pipe_in_en                (pipein_en),
        .pipe_out_data             (pipeout),      
        .pipe_out_read             (pipeout_en),
        .cfg                       (cfg),
        .data_stream_en            (stream_en),
        .status                    (status)                
        );

    always #1 clk=~clk;
 
 
     initial begin
        #16     pipein_en  = 1;
                pipein     = 16'h0200;
        
        #2      pipein     = 16'h1234;
        
        #2      pipein     = 16'h0100;
        
        #2      pipein     = 16'h0101;
        
        #2      pipein     = 16'h0102;  // should read 'no error' (0)
        
        #2      pipein     = 16'h0100;
        
        #2      pipein     = 16'h0101;
                
        #2      pipein     = 16'h01F1;
                
        #2      pipein     = 16'h0102; // should read 'unknown command' (1)

        #2      pipein     = 16'h0102; // should read 'no error' (0)

        #2      pipein     = 16'h0101;

        #2      pipein     = 16'h0100;

        #2      pipein     = 16'h0101;

        #2      pipein     = 16'h0101;

        #2      pipein_en  = 0;
        
        #2      pipeout_en = 1;
        
        #2      pipeout_en = 0;
        
        #4      pipeout_en = 1;
        
        #6      pipeout_en = 0;
         
        #2      pipein_en  = 1;
                pipein     = 16'h0102;  // should read 'FIFO full' (2)

        #2      pipein_en  = 0;
        
        #4      pipeout_en = 1;
        
        #20     pipein_en  = 1;
                pipein     = 16'h0102;  // should read 'FIFO empty' (4)

        #2      pipein_en  = 0;
         
    end
 
 
 
 
 
    initial begin
                reset      = 0;

        #4      reset      = 1;
        
        #2      reset      = 0;
                stream_en  = 8'h12;
                pipein     = 16'h0000;
                pipein_en  = 0;
                pipeout_en = 0;
                cfg        = 16'h0000;
        
        #4      data_write    = 1;
                data_to_write = header_magic_number[15:0];
        
        #2      data_to_write = header_magic_number[31:16];
        
        #2      data_to_write = header_magic_number[47:32];
        
        #2      data_to_write = header_magic_number[63:48];
        
        #2      data_to_write = 16'h4401;    // timestamp
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4402;
                data_write    = 1;
        #2      data_write    = 0;


        #2      data_to_write = 16'h4200;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4201;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4202;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4203;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4204;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4205;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4206;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4207;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4208;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4209;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h420A;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h420B;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h420C;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h420D;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h420E;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h420F;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4210;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4211;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4212;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4213;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4214;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4215;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4216;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4217;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4218;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4219;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h421A;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h421B;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h421C;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h421D;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h421E;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h421F;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4220;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4221;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4222;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4223;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4224;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4225;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4226;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4227;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4228;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4229;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h422A;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h422B;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h422C;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h422D;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h422E;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h422F;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4230;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4231;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4232;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4233;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4234;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4235;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4236;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4237;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4238;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4239;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h423A;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h423B;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h423C;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h423D;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h423E;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h423F;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4240;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4241;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4242;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4243;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4244;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4245;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4246;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4247;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4248;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4249;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h424A;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h424B;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h424C;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h424D;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h424E;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h424F;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4250;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4251;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4252;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4254;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4253;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4255;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4256;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4257;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4258;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h4259;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h425A;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h425B;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h425C;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h425D;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h425E;
                data_write    = 1;
        #2      data_write    = 0;

        #2      data_to_write = 16'h425F;
        #2      data_to_write = 16'h4260;
        #2      data_to_write = 16'h4261;
        #2      data_to_write = 16'h4262;
        #2      data_to_write = 16'h4263;
        #2      data_to_write = 16'h4264;
        #2      data_to_write = 16'h4265;
        #2      data_to_write = 16'h4266;
        #2      data_to_write = 16'h4267;
        #2      data_to_write = 16'h4268;
        #2      data_to_write = 16'h4269;
        #2      data_to_write = 16'h426A;
        #2      data_to_write = 16'h426B;
        #2      data_to_write = 16'h426C;
        #2      data_to_write = 16'h426D;
        #2      data_to_write = 16'h426E;
        #2      data_to_write = 16'h426F;
        #2      data_to_write = 16'h4270;
        #2      data_to_write = 16'h4271;
        #2      data_to_write = 16'h4272;
        #2      data_to_write = 16'h4273;
        #2      data_to_write = 16'h4274;
        #2      data_to_write = 16'h4275;
        #2      data_to_write = 16'h4276;
        #2      data_to_write = 16'h4277;
        #2      data_to_write = 16'h4278;
        #2      data_to_write = 16'h4279;
        #2      data_to_write = 16'h427A;
        #2      data_to_write = 16'h427B;
        #2      data_to_write = 16'h427C;
        #2      data_to_write = 16'h427D;
        #2      data_to_write = 16'h427E;
        #2      data_to_write = 16'h427F;
        #2      data_to_write = 16'h4280;
        #2      data_to_write = 16'h4281;
        #2      data_to_write = 16'h4282;
        #2      data_to_write = 16'h4283;
        #2      data_to_write = 16'h4284;
        #2      data_to_write = 16'h4285;
        #2      data_to_write = 16'h4286;
        #2      data_to_write = 16'h4287;
        #2      data_to_write = 16'h4288;
        #2      data_to_write = 16'h4289;
        #2      data_to_write = 16'h428A;
        #2      data_to_write = 16'h428B;
        #2      data_to_write = 16'h428C;
        #2      data_to_write = 16'h428D;
        #2      data_to_write = 16'h428E;
        #2      data_to_write = 16'h428F;
        #2      data_to_write = 16'h4290;
        #2      data_to_write = 16'h4291;
        #2      data_to_write = 16'h4292;
        #2      data_to_write = 16'h4293;
        #2      data_to_write = 16'h4294;
        #2      data_to_write = 16'h4295;
        #2      data_to_write = 16'h4296;
        #2      data_to_write = 16'h4297;
        #2      data_to_write = 16'h4298;
        #2      data_to_write = 16'h4299;
        #2      data_to_write = 16'h429A;
        #2      data_to_write = 16'h429B;
        #2      data_to_write = 16'h429C;
        #2      data_to_write = 16'h429D;
        #2      data_to_write = 16'h429E;
        #2      data_to_write = 16'h429F;
        #2      data_to_write = 16'h42A0;
        #2      data_to_write = 16'h42A1;
        #2      data_to_write = 16'h42A2;
        #2      data_to_write = 16'h42A3;
        #2      data_to_write = 16'h42A4;
        #2      data_to_write = 16'h42A5;
        #2      data_to_write = 16'h42A6;
        #2      data_to_write = 16'h42A7;
        #2      data_to_write = 16'h42A8;
        #2      data_to_write = 16'h42A9;
        #2      data_to_write = 16'h42AA;
        #2      data_to_write = 16'h42AB;
        #2      data_to_write = 16'h42AC;
        #2      data_to_write = 16'h42AD;
        #2      data_to_write = 16'h42AE;
        #2      data_to_write = 16'h42AF;
        #2      data_to_write = 16'h42B0;
        #2      data_to_write = 16'h42B1;
        #2      data_to_write = 16'h42B2;
        #2      data_to_write = 16'h42B3;
        #2      data_to_write = 16'h42B4;
        #2      data_to_write = 16'h42B5;
        #2      data_to_write = 16'h42B6;
        #2      data_to_write = 16'h42B7;
        #2      data_to_write = 16'h42B8;
        #2      data_to_write = 16'h42B9;
        #2      data_to_write = 16'h42BA;
        #2      data_to_write = 16'h42BB;
        #2      data_to_write = 16'h42BC;
        #2      data_to_write = 16'h42BD;
        #2      data_to_write = 16'h42BE;
        #2      data_to_write = 16'h42BF;
        #2      data_to_write = 16'h42C0;
        #2      data_to_write = 16'h42C1;
        #2      data_to_write = 16'h42C2;
        #2      data_to_write = 16'h42C3;
        #2      data_to_write = 16'h42C4;
        #2      data_to_write = 16'h42C5;
        #2      data_to_write = 16'h42C6;
        #2      data_to_write = 16'h42C7;
        #2      data_to_write = 16'h42C8;
        #2      data_to_write = 16'h42C9;
        #2      data_to_write = 16'h42CA;
        #2      data_to_write = 16'h42CB;
        #2      data_to_write = 16'h42CC;
        #2      data_to_write = 16'h42CD;
        #2      data_to_write = 16'h42CE;
        #2      data_to_write = 16'h42CF;
        #2      data_to_write = 16'h42D0;
        #2      data_to_write = 16'h42D1;
        #2      data_to_write = 16'h42D2;
        #2      data_to_write = 16'h42D3;
        #2      data_to_write = 16'h42D4;
        #2      data_to_write = 16'h42D5;
        #2      data_to_write = 16'h42D6;
        #2      data_to_write = 16'h42D7;
        #2      data_to_write = 16'h42D8;
        #2      data_to_write = 16'h42D9;
        #2      data_to_write = 16'h42DA;
        #2      data_to_write = 16'h42DB;
        #2      data_to_write = 16'h42DC;
        #2      data_to_write = 16'h42DD;
        #2      data_to_write = 16'h42DE;
        #2      data_to_write = 16'h42DF;
        #2      data_to_write = 16'h42E0;
        #2      data_to_write = 16'h42E1;
        #2      data_to_write = 16'h42E2;
        #2      data_to_write = 16'h42E3;
        #2      data_to_write = 16'h42E4;
        #2      data_to_write = 16'h42E5;
        #2      data_to_write = 16'h42E6;
        #2      data_to_write = 16'h42E7;
        #2      data_to_write = 16'h42E8;
        #2      data_to_write = 16'h42E9;
        #2      data_to_write = 16'h42EA;
        #2      data_to_write = 16'h42EB;
        #2      data_to_write = 16'h42EC;
        #2      data_to_write = 16'h42ED;
        #2      data_to_write = 16'h42EE;
        #2      data_to_write = 16'h42EF;
        #2      data_to_write = 16'h42F0;
        #2      data_to_write = 16'h42F1;
        #2      data_to_write = 16'h42F2;
        #2      data_to_write = 16'h42F3;
        #2      data_to_write = 16'h42F4;
        #2      data_to_write = 16'h42F5;
        #2      data_to_write = 16'h42F6;
        #2      data_to_write = 16'h42F7;
        #2      data_to_write = 16'h42F8;
        #2      data_to_write = 16'h42F9;
        #2      data_to_write = 16'h42FA;
        #2      data_to_write = 16'h42FB;
        #2      data_to_write = 16'h42FC;
        #2      data_to_write = 16'h42FD;
        #2      data_to_write = 16'h42FE;
        #2      data_to_write = 16'h42FF;
        #2      data_to_write = 16'h6900;
        #2      data_to_write = 16'h6901;
        #2      data_to_write = 16'h6902;
        #2      data_to_write = 16'h6903;
        #2      data_to_write = 16'h6904;
        #2      data_to_write = 16'h6905;
        #2      data_to_write = 16'h6906;
        #2      data_to_write = 16'h6907;
        #2      data_to_write = 16'h6908;
        #2      data_to_write = 16'h6909;
        #2      data_to_write = 16'h690A;
        #2      data_to_write = 16'h690B;
        #2      data_to_write = 16'h690C;
        #2      data_to_write = 16'h690D;
        #2      data_to_write = 16'h690E;
        #2      data_to_write = 16'h690F;
        #2      data_to_write = 16'h6910;
        #2      data_to_write = 16'h6911;
        #2      data_to_write = 16'h6912;
        #2      data_to_write = 16'h6913;
        #2      data_to_write = 16'h6914;
        #2      data_to_write = 16'h6915;
        #2      data_to_write = 16'h6916;
        #2      data_to_write = 16'h6917;
        #2      data_to_write = 16'h6918;
        #2      data_to_write = 16'h6919;
        #2      data_to_write = 16'h691A;
        #2      data_to_write = 16'h691B;
        #2      data_to_write = 16'h691C;
        #2      data_to_write = 16'h691D;
        #2      data_to_write = 16'h691E;
        #2      data_to_write = 16'h691F;
        #2      data_to_write = 16'h6920;
        #2      data_to_write = 16'h6921;
        #2      data_to_write = 16'h6922;
        #2      data_to_write = 16'h6923;
        #2      data_to_write = 16'h6924;
        #2      data_to_write = 16'h6925;
        #2      data_to_write = 16'h6926;
        #2      data_to_write = 16'h6927;
        #2      data_to_write = 16'h6928;
        #2      data_to_write = 16'h6929;
        #2      data_to_write = 16'h692A;
        #2      data_to_write = 16'h692B;
        #2      data_to_write = 16'h692C;
        #2      data_to_write = 16'h692D;
        #2      data_to_write = 16'h692E;
        #2      data_to_write = 16'h692F;
        #2      data_to_write = 16'h6930;
        #2      data_to_write = 16'h6931;
        #2      data_to_write = 16'h6932;
        #2      data_to_write = 16'h6933;
        #2      data_to_write = 16'h6934;
        #2      data_to_write = 16'h6935;
        #2      data_to_write = 16'h6936;
        #2      data_to_write = 16'h6937;
        #2      data_to_write = 16'h6938;
        #2      data_to_write = 16'h6939;
        #2      data_to_write = 16'h693A;
        #2      data_to_write = 16'h693B;
        #2      data_to_write = 16'h693C;
        #2      data_to_write = 16'h693D;
        #2      data_to_write = 16'h693E;
        #2      data_to_write = 16'h693F;
        #2      data_to_write = 16'h6940;
        #2      data_to_write = 16'h6941;
        #2      data_to_write = 16'h6942;
        #2      data_to_write = 16'h6943;
        #2      data_to_write = 16'h6944;
        #2      data_to_write = 16'h6945;
        #2      data_to_write = 16'h6946;
        #2      data_to_write = 16'h6947;
        #2      data_to_write = 16'h6948;
        #2      data_to_write = 16'h6949;
        #2      data_to_write = 16'h694A;
        #2      data_to_write = 16'h694B;
        #2      data_to_write = 16'h694C;
        #2      data_to_write = 16'h694D;
        #2      data_to_write = 16'h694E;
        #2      data_to_write = 16'h694F;
        #2      data_to_write = 16'h6950;
        #2      data_to_write = 16'h6951;
        #2      data_to_write = 16'h6952;
        #2      data_to_write = 16'h6953;
        #2      data_to_write = 16'h6954;
        #2      data_to_write = 16'h6955;
        #2      data_to_write = 16'h6956;
        #2      data_to_write = 16'h6957;
        #2      data_to_write = 16'h6958;
        #2      data_to_write = 16'h6959;
        #2      data_to_write = 16'h695A;
        #2      data_to_write = 16'h695B;
        #2      data_to_write = 16'h695C;
        #2      data_to_write = 16'h695D;
        #2      data_to_write = 16'h695E;
        #2      data_to_write = 16'h695F;
        #2      data_to_write = 16'h6960;
        #2      data_to_write = 16'h6961;
        #2      data_to_write = 16'h6962;
        #2      data_to_write = 16'h6963;
        #2      data_to_write = 16'h6964;
        #2      data_to_write = 16'h6965;
        #2      data_to_write = 16'h6966;
        #2      data_to_write = 16'h6967;
        #2      data_to_write = 16'h6968;
        #2      data_to_write = 16'h6969;
        #2      data_to_write = 16'h696A;
        #2      data_to_write = 16'h696B;
        #2      data_to_write = 16'h696C;
        #2      data_to_write = 16'h696D;
        #2      data_to_write = 16'h696E;
        #2      data_to_write = 16'h696F;
        #2      data_to_write = 16'h6970;
        #2      data_to_write = 16'h6971;
        #2      data_to_write = 16'h6972;
        #2      data_to_write = 16'h6973;
        #2      data_to_write = 16'h6974;
        #2      data_to_write = 16'h6975;
        #2      data_to_write = 16'h6976;
        #2      data_to_write = 16'h6977;
        #2      data_to_write = 16'h6978;
        #2      data_to_write = 16'h6979;
        #2      data_to_write = 16'h697A;
        #2      data_to_write = 16'h697B;
        #2      data_to_write = 16'h697C;
        #2      data_to_write = 16'h697D;
        #2      data_to_write = 16'h697E;
        #2      data_to_write = 16'h697F;
        #2      data_to_write = 16'h6980;
        #2      data_to_write = 16'h6981;
        #2      data_to_write = 16'h6982;
        #2      data_to_write = 16'h6983;
        #2      data_to_write = 16'h6984;
        #2      data_to_write = 16'h6985;
        #2      data_to_write = 16'h6986;
        #2      data_to_write = 16'h6987;
        #2      data_to_write = 16'h6988;
        #2      data_to_write = 16'h6989;
        #2      data_to_write = 16'h698A;
        #2      data_to_write = 16'h698B;
        #2      data_to_write = 16'h698C;
        #2      data_to_write = 16'h698D;
        #2      data_to_write = 16'h698E;
        #2      data_to_write = 16'h698F;
        #2      data_to_write = 16'h6990;
        #2      data_to_write = 16'h6991;
        #2      data_to_write = 16'h6992;
        #2      data_to_write = 16'h6993;
        #2      data_to_write = 16'h6994;
        #2      data_to_write = 16'h6995;
        #2      data_to_write = 16'h6996;
        #2      data_to_write = 16'h6997;
        #2      data_to_write = 16'h6998;
        #2      data_to_write = 16'h6999;
        #2      data_to_write = 16'h699A;
        #2      data_to_write = 16'h699B;
        #2      data_to_write = 16'h699C;
        #2      data_to_write = 16'h699D;
        #2      data_to_write = 16'h699E;
        #2      data_to_write = 16'h699F;
        #2      data_to_write = 16'h69A0;
        #2      data_to_write = 16'h69A1;
        #2      data_to_write = 16'h69A2;
        #2      data_to_write = 16'h69A3;
        #2      data_to_write = 16'h69A4;
        #2      data_to_write = 16'h69A5;
        #2      data_to_write = 16'h69A6;
        #2      data_to_write = 16'h69A7;
        #2      data_to_write = 16'h69A8;
        #2      data_to_write = 16'h69A9;
        #2      data_to_write = 16'h69AA;
        #2      data_to_write = 16'h69AB;
        #2      data_to_write = 16'h69AC;
        #2      data_to_write = 16'h69AD;
        #2      data_to_write = 16'h69AE;
        #2      data_to_write = 16'h69AF;
        #2      data_to_write = 16'h69B0;
        #2      data_to_write = 16'h69B1;
        #2      data_to_write = 16'h69B2;
        #2      data_to_write = 16'h69B3;
        #2      data_to_write = 16'h69B4;
        #2      data_to_write = 16'h69B5;
        #2      data_to_write = 16'h69B6;
        #2      data_to_write = 16'h69B7;
        #2      data_to_write = 16'h69B8;
        #2      data_to_write = 16'h69B9;
        #2      data_to_write = 16'h69BA;
        #2      data_to_write = 16'h69BB;
        #2      data_to_write = 16'h69BC;
        #2      data_to_write = 16'h69BD;
        #2      data_to_write = 16'h69BE;
        #2      data_to_write = 16'h69BF;
        #2      data_to_write = 16'h69C0;
        #2      data_to_write = 16'h69C1;
        #2      data_to_write = 16'h69C2;
        #2      data_to_write = 16'h69C3;
        #2      data_to_write = 16'h69C4;
        #2      data_to_write = 16'h69C5;
        #2      data_to_write = 16'h69C6;
        #2      data_to_write = 16'h69C7;
        #2      data_to_write = 16'h69C8;
        #2      data_to_write = 16'h69C9;
        #2      data_to_write = 16'h69CA;
        #2      data_to_write = 16'h69CB;
        #2      data_to_write = 16'h69CC;
        #2      data_to_write = 16'h69CD;
        #2      data_to_write = 16'h69CE;
        #2      data_to_write = 16'h69CF;
        #2      data_to_write = 16'h69D0;
        #2      data_to_write = 16'h69D1;
        #2      data_to_write = 16'h69D2;
        #2      data_to_write = 16'h69D3;
        #2      data_to_write = 16'h69D4;
        #2      data_to_write = 16'h69D5;
        #2      data_to_write = 16'h69D6;
        #2      data_to_write = 16'h69D7;
        #2      data_to_write = 16'h69D8;
        #2      data_to_write = 16'h69D9;
        #2      data_to_write = 16'h69DA;
        #2      data_to_write = 16'h69DB;
        #2      data_to_write = 16'h69DC;
        #2      data_to_write = 16'h69DD;
        #2      data_to_write = 16'h69DE;
        #2      data_to_write = 16'h69DF;
        #2      data_to_write = 16'h69E0;
        #2      data_to_write = 16'h69E1;
        #2      data_to_write = 16'h69E2;
        #2      data_to_write = 16'h69E3;
        #2      data_to_write = 16'h69E4;
        #2      data_to_write = 16'h69E5;
        #2      data_to_write = 16'h69E6;
        #2      data_to_write = 16'h69E7;
        #2      data_to_write = 16'h69E8;
        #2      data_to_write = 16'h69E9;
        #2      data_to_write = 16'h69EA;
        #2      data_to_write = 16'h69EB;
        #2      data_to_write = 16'h69EC;
        #2      data_to_write = 16'h69ED;
        #2      data_to_write = 16'h69EE;
        #2      data_to_write = 16'h69EF;
        #2      data_to_write = 16'h69F0;
        #2      data_to_write = 16'h69F1;
        #2      data_to_write = 16'h69F2;
        #2      data_to_write = 16'h69F3;
        #2      data_to_write = 16'h69F4;
        #2      data_to_write = 16'h69F5;
        #2      data_to_write = 16'h69F6;
        #2      data_to_write = 16'h69F7;
        #2      data_to_write = 16'h69F8;
        #2      data_to_write = 16'h69F9;
        #2      data_to_write = 16'h69FA;
        #2      data_to_write = 16'h69FB;
        #2      data_to_write = 16'h69FC;
        #2      data_to_write = 16'h69FD;
        #2      data_to_write = 16'h69FE;
        #2      data_to_write = 16'h69FF;
        $finish;
    end
 
endmodule